module zero
(
output [15:0] out
);

assign out[15:0] = 0;

endmodule