module decoder
(

	input A,
	output B
);

assign B = A;
endmodule